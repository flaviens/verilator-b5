module top(in_data, out_data);
  wire _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire [209:0] _086_;
  wire [131:0] _087_;
  wire [131:0] _088_;
  wire [234:0] _089_;
  wire [234:0] _090_;
  wire [234:0] _091_;
  wire [52:0] _092_;
  wire [47:0] _093_;
  wire [74:0] _094_;
  wire [74:0] _095_;
  wire [74:0] _096_;
  wire [47:0] _097_;
  wire [90:0] _098_;
  wire [90:0] _099_;
  wire [269:0] _100_;
  wire [269:0] _101_;
  wire [51:0] _102_;
  wire [228:0] _103_;
  wire [228:0] _104_;
  wire [228:0] _105_;
  wire [170:0] _106_;
  wire [170:0] _107_;
  wire [23:0] _108_;
  wire [23:0] _109_;
  wire [162:0] _110_;
  wire [276:0] _111_;
  wire [276:0] _112_;
  wire [227:0] _113_;
  wire [60:0] _114_;
  wire [60:0] _115_;
  wire [152:0] _116_;
  wire [228:0] _117_;
  wire [282:0] _118_;
  wire [282:0] _119_;
  wire [264:0] _120_;
  wire [217:0] _121_;
  wire [260:0] _122_;
  wire [260:0] _123_;
  wire [267:0] _124_;
  wire [148:0] _125_;
  wire [22:0] _126_;
  wire [295:0] _127_;
  wire [206:0] _128_;
  wire [91:0] _129_;
  wire [164:0] _130_;
  wire [100:0] _131_;
  wire [210:0] _132_;
  wire [170:0] _133_;
  wire [210:0] _134_;
  wire [222:0] _135_;
  wire [288:0] _136_;
  wire [161:0] _137_;
  wire [161:0] _138_;
  wire [59:0] _139_;
  wire [59:0] _140_;
  wire [278:0] _141_;
  wire [278:0] _142_;
  wire [210:0] _143_;
  wire [21:0] _144_;
  wire [286:0] _145_;
  wire [211:0] _146_;
  input [2399:0] in_data;
  wire [2399:0] in_data;
  output [895:0] out_data;
  wire [895:0] out_data;
  assign _000_ = _002_ ^ _001_;
  assign _003_ = _005_ ^ _004_;
  assign _006_ = _008_ ^ _007_;
  assign _009_ = _010_ ^ _006_;
  assign _011_ = _013_ ^ _012_;
  assign _014_ = _016_ ^ _015_;
  assign _017_ = _019_ ^ _018_;
  assign _020_ = _022_ ^ _021_;
  assign _023_ = _011_ ^ _024_;
  assign _025_ = _026_ ^ _011_;
  assign _027_ = _029_ ^ _028_;
  assign _030_ = in_data[110] ^ _031_;
  assign _004_ = _012_ ^ _032_;
  assign _033_ = _000_ ^ _004_;
  assign _034_ = _036_ ^ _035_;
  assign _037_ = _027_ ^ _038_;
  assign _039_ = _041_ ^ _040_;
  assign _042_ = _044_ ^ _043_;
  assign _045_ = _047_ ^ _046_;
  assign _048_ = _033_ ^ _002_;
  assign _049_ = _050_ ^ _020_;
  assign _051_ = _009_ ^ _025_;
  assign _052_ = _053_ ^ _012_;
  assign _054_ = _022_ ^ _055_;
  assign _056_ = _006_ ^ _057_;
  assign out_data[832] = _049_ ^ _059_;
  assign out_data[768] = _024_ ^ _060_;
  assign out_data[736] = _020_ ^ _062_;
  assign out_data[672] = _064_ ^ in_data[381];
  assign _058_ = _063_ ^ _061_;
  assign out_data[576] = _066_ ^ _065_;
  assign out_data[544] = _030_ ^ out_data[672];
  assign out_data[480] = _068_ ^ _067_;
  assign out_data[416] = _039_ ^ _023_;
  assign out_data[320] = _058_ ^ _045_;
  assign out_data[256] = _037_ ^ _069_;
  assign out_data[224] = _034_ ^ _070_;
  assign out_data[96] = in_data[2290] ^ _072_;
  assign out_data[64] = _073_ ^ out_data[224];
  assign out_data[32] = _076_ ^ _075_;
  assign out_data[0] = _077_ ^ _000_;
  assign _069_ = _074_ ^ _071_;
  assign _022_ = _078_ ^ _069_;
  assign _079_ = _081_ ^ _080_;
  assign _055_ = _082_ ^ _069_;
  assign _012_ = in_data[1512] ^ in_data[117];
  assign _083_ = _079_ ^ _055_;
  assign _024_ = _084_ ^ _012_;
  assign _036_ = _085_ ^ _055_;
  assign { _123_[125:109], _104_[228:136], _123_[15:0] } = { _112_[244:216], _095_[74:2], _005_, _117_[24:2] } + { _088_[109:45], _019_, _088_[43:1], _107_[16:3], _024_, _004_, _055_ };
  assign { _087_[131:123], _035_, _087_[121:0] } = { _086_[180:89], _032_, _086_[87:49] } + { _088_[131:45], _019_, _088_[43:1], _036_ };
  assign { _089_[234:161], _018_, _089_[159:123], _015_, _089_[121:0] } = { _091_[234:198], _087_[131:123], _035_, _087_[121:0], _091_[65:58], _016_, _091_[56:43], _085_, _091_[41:32], _062_, _091_[30:23], _007_, _091_[21:1], _003_ } + { _086_[89], _032_, _086_[87:40], _074_, _086_[38:30], _090_[174:105], _066_, _090_[103:40], _004_, _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0] };
  assign { _134_[155:131], _097_[47], _001_, _097_[45:22], _096_[74:39], _063_, _096_[37:6], _134_[35:23], _010_, _134_[21:1] } = { in_data[720:567], _012_ } + in_data[1712:1558];
  assign { _092_[52:35], _068_, _092_[33:17], _028_, _092_[15:0] } = { _087_[107:56], _058_ } + { _087_[118:67], _012_ };
  assign { _094_[74:14], _046_, _026_, _094_[11:0] } = { _096_[74:39], _063_, _096_[37:6], _079_, _022_, _003_, _058_, _055_, _022_ } + _095_;
  assign { _098_[90:58], _029_, _098_[56:0] } = { _089_[114:26], _009_, _055_ } + { _095_[63:0], _099_[26:4], _059_, _099_[2:0] };
  assign { _100_[269:129], _057_, _100_[127:0] } = { _101_[269:169], _076_, _101_[167:158], _091_[234:218], _098_[90:58], _029_, _098_[56:0], _058_, _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _079_ } + { _098_[84:58], _029_, _098_[56:28], _079_, _086_[209:89], _032_, _086_[87:40], _074_, _086_[38:0], _083_, _058_ };
  assign { _102_[51:33], _021_, _102_[31:0] } = _101_[251:200] + { _091_[65:58], _016_, _091_[56:43], _085_, _091_[41:32], _062_, _091_[30:23], _007_, _091_[21:14] };
  assign { _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0] } = { in_data[1326:1280], _012_ } + { _097_[47], _001_, _097_[45:22], _096_[74:53] };
  assign _103_ = { _101_[202:169], _076_, _101_[167:158], _091_[234:204], _091_[65:58], _016_, _091_[56:43], _085_, _091_[41:32], _062_, _091_[30:23], _007_, _091_[21:1], _020_, _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_, _094_[74:14], _046_, _026_, _094_[11:0] } + { _104_[228:136], _083_, _036_, _087_[131:123], _035_, _087_[121:0], _009_, _036_ };
  assign { _106_[170:42], _065_, _106_[40:0] } = { _107_[170:148], _088_[131:45], _019_, _088_[43:1], _107_[16:1], _014_ } + { _090_[168:158], _079_, _055_, _027_, _020_, _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _009_, _020_, _092_[52:35], _068_, _092_[33:17], _028_, _092_[15:0], _092_[52:35], _068_, _092_[33:17], _028_, _092_[15:0] };
  assign { _108_[23], _041_, _108_[21:20], _043_, _108_[18:0] } = { _088_[47:45], _019_, _088_[43:25], _009_ } + { _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4], _069_, _055_, _003_, _022_ };
  assign { _047_, _110_[161:0] } = { _101_[204:169], _076_, _101_[167:158], _091_[234:211], _102_[51:33], _021_, _102_[31:0], _027_, _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0] } + { _106_[59:42], _065_, _106_[40:1], _009_, _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0], _102_[51:33], _021_, _102_[31:0], _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_ };
  assign _111_ = { _103_[227:53], _036_, _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _092_[52:35], _068_, _092_[33:17], _028_, _092_[15:0] } + { _112_[276:216], _095_, _099_[26:22], _090_[174:105], _066_, _090_[103:40], _000_ };
  assign _113_ = { _095_[35:0], _099_[26:6], _106_[170:42], _065_, _106_[40:0] } + { _091_[64:58], _016_, _091_[56:52], _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0], _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0], _090_[174:105], _066_, _090_[103:40], _020_, _027_ };
  assign _114_ = { _115_[60:6], _031_, _115_[4:2], _069_, _011_ } + { _090_[139:105], _066_, _090_[103:79] };
  assign { _116_[152:37], _050_, _116_[35:15], _073_, _116_[13:0] } = in_data[740:588] + { _087_[64:62], _094_[74:14], _046_, _026_, _094_[11:0], _094_[74:14], _046_, _026_, _094_[11:0] };
  assign { _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_ } = { _086_[195:185], _004_ } + _086_[189:178];
  assign _118_ = { _119_[282:255], _081_, _119_[253:25], _108_[23], _041_, _108_[21:20], _043_, _108_[18:0], _058_ } + { _113_[184:158], _103_, _025_, _108_[23], _041_, _108_[21:20], _043_, _108_[18:0], _083_, _004_ };
  assign { _121_[217:73], _064_, _121_[71:0] } = _113_[219:2] + { _086_[185:89], _032_, _086_[87:40], _074_, _086_[38:32], _048_, _014_, _114_, _049_ };
  assign _122_ = { _120_[259:258], _119_[282:255], _081_, _119_[253:25], _017_ } + { _115_[38:6], _031_, _115_[4:2], _123_[223:129], _051_, _045_, _052_, _123_[125:109], _104_[228:136], _123_[15:0] };
  assign { _120_[264:258], _119_[282:255], _081_, _119_[253:25] } = { in_data[1705:1651], _086_[209:89], _032_, _086_[87:40], _074_, _086_[38:0] } + in_data[2254:1990];
  assign _125_ = { _106_[133:42], _065_, _106_[40:9], _108_[23], _041_, _108_[21:20], _043_, _108_[18:0] } + { _111_[156:9], _079_ };
  assign _126_ = { _092_[32:17], _028_, _092_[15:10] } + { _092_[48:35], _068_, _092_[33:26] };
  assign { _127_[295:220], out_data[831:800], _127_[187:157], _060_, _127_[155], _067_, _127_[153:0] } = { _088_[100:91], _042_, _052_, _118_, _051_ } + { _111_[140:85], _045_, _102_[51:33], _021_, _102_[31:0], _047_, _110_[161:0], _126_, _027_ };
  assign { _128_[206:203], out_data[735:704], _128_[170:0] } = { _113_[218:64], _102_[51:33], _021_, _102_[31:0] } + { in_data[860:793], _055_, _094_[74:14], _046_, _026_, _094_[11:0], _114_, _030_, _058_ };
  assign { _129_[91:44], out_data[671:640], _129_[11:0] } = _122_[109:18] + { _116_[103:37], _050_, _116_[35:15], _073_, _116_[13:12] };
  assign { _130_[164:136], out_data[639:608], _130_[103:31], _072_, _130_[29:0] } = { _104_[195:190], _090_[174:105], _066_, _090_[103:40], _108_[23], _041_, _108_[21:20], _043_, _108_[18:0] } + _122_[252:88];
  assign { _131_[100:92], _077_, _131_[90:82], out_data[543:512], _131_[49:0] } = { _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _012_, _102_[51:33], _021_, _102_[31:0] } + { _123_[110:109], _104_[228:136], _123_[15:11], out_data[736] };
  assign { _133_[170:125], out_data[479:448], _133_[92:59], _075_, _133_[57:0] } = { _106_[170:42], _065_, _106_[40:0] } + { _089_[181:161], _018_, _089_[159:123], _015_, _089_[121:11] };
  assign { _135_[222:181], out_data[415:384], _135_[148:71], _070_, _135_[69:0] } = { _123_[124:109], _104_[228:136], _123_[15:1], _108_[23], _041_, _108_[21:20], _043_, _108_[18:0], _091_[65:58], _016_, _091_[56:43], _085_, _091_[41:32], _062_, _091_[30:23], _007_, _091_[21:1], _004_, _052_, out_data[672], _054_, _036_, _023_, _054_, _023_, out_data[832], out_data[416] } + { _110_[148:21], _034_, _129_[91:44], out_data[671:640], _129_[11:0], _052_, out_data[416] };
  assign { _136_[288:225], out_data[383:352], _136_[192:0] } = { in_data[2157:2076], _128_[206:203], out_data[735:704], _128_[170:0] } + { _128_[166:30], _012_, _025_, _055_, _125_ };
  assign { _132_[210], _084_, _132_[208:159], _115_[60:6], _031_, _115_[4:2], _123_[223:129], _132_[4:0] } = { in_data[1114:917], _004_, _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_ } + { _093_[13:10], _058_, _012_, _058_, _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _134_[155:131], _097_[47], _001_, _097_[45:22], _096_[74:39], _063_, _096_[37:6], _134_[35:23], _010_, _134_[21:1], _012_ };
  assign { _137_[161:39], out_data[319:288], _137_[6:0] } = { _118_[162:2], out_data[832] } + { _095_[39:0], _099_[26:4], _059_, _099_[2:0], _124_[128:92], _138_[57:49], _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], out_data[320] };
  assign { _139_[59:49], out_data[223:192], _139_[16:0] } = { _140_[59:47], _101_[269:224], _045_ } + { _101_[204:171], _017_, _052_, _005_, _117_[24:2] };
  assign { _141_[278:37], out_data[191:160], _141_[4:0] } = { _087_[126:123], _035_, _087_[121:102], _142_[253:247], _107_[170:148], _088_[131:45], _019_, _088_[43:1], _107_[16:1], _142_[76:0] } + { _103_[215:16], _094_[74:14], _046_, _026_, _094_[11:0], _049_, _056_, _051_, out_data[544] };
  assign { _143_[210:163], out_data[159:128], _143_[130:0] } = { _086_[191:89], _032_, _086_[87:40], _074_, _086_[38:19], _036_, _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_, _005_, _117_[24:2], _012_ } + { _118_[255:47], out_data[576], out_data[544] };
  assign { _086_[209:89], _032_, _086_[87:40], _074_, _086_[38:0] } = in_data[801:592] + in_data[1802:1593];
  assign { _040_, _144_[20], _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4] } = { in_data[2200:2180], _069_ } + in_data[711:690];
  assign { _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0] } = { _097_[24:22], _096_[74:40], _004_ } + { _093_[30:9], _082_, _093_[7:6], _069_, _004_, _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_ };
  assign { _090_[174:105], _066_, _090_[103:40] } = { _086_[117:89], _032_, _086_[87:40], _074_, _086_[38:6], _040_, _144_[20], _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4], _058_ } + { _132_[190:159], _115_[60:6], _031_, _115_[4:2], _123_[223:204], _079_, _040_, _144_[20], _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4], _012_ };
  assign { _145_[286:250], _112_[276:216], _095_, _099_[26:4], _059_, _099_[2:0], _124_[128:92], _138_[57:49], _145_[40:0] } = { in_data[1464:1262], _055_, _012_, _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0], _022_, _012_, _058_, _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0], _079_ } + { _115_[45:6], _031_, _115_[4:2], _123_[223:136], _134_[155:131], _097_[47], _001_, _097_[45:22], _096_[74:39], _063_, _096_[37:6], _134_[35:23], _010_, _134_[21:1] };
  assign { _091_[65:58], _016_, _091_[56:43], _085_, _091_[41:32], _062_, _091_[30:23], _007_, _091_[21:1] } = { _145_[263:250], _112_[276:227], _012_ } + { _090_[142:105], _066_, _090_[103:78] };
  assign { _146_[211:189], _140_[59:47], _101_[269:169], _076_, _101_[167:158], _091_[234:198], _146_[26:0] } = { _119_[239:50], _040_, _144_[20], _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4] } + { _119_[237:27], _058_ };
  assign { _142_[253:247], _107_[170:148], _088_[131:45], _019_, _088_[43:1], _107_[16:1], _142_[76:0] } = { _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _132_[210], _084_, _132_[208:159], _115_[60:6], _031_, _115_[4:2], _123_[223:129], _132_[4:0], _058_ } + { _086_[83:40], _074_, _086_[38:36], _004_, _055_, _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_, _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_, _022_, _055_, _079_, _040_, _144_[20], _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4], _134_[155:131], _097_[47], _001_, _097_[45:22], _096_[74:39], _063_, _096_[37:6], _134_[35:23], _010_, _134_[21:1] };
  assign { _005_, _117_[24:2] } = { _091_[30:23], _007_, _091_[21:7] } + { _090_[63:52], _105_[86:84], _044_, _105_[82:79], _071_, _105_[77:76], _078_ };
  assign { _086_[88], _086_[39] } = { _032_, _074_ };
  assign _087_[122] = _035_;
  assign { _088_[44], _088_[0] } = { _019_, _036_ };
  assign { _089_[160], _089_[122] } = { _018_, _015_ };
  assign { _090_[234:175], _090_[104], _090_[39], _090_[29], _090_[8] } = { _086_[89], _032_, _086_[87:40], _074_, _086_[38:30], _066_, _004_, _008_, _002_ };
  assign { _091_[197:66], _091_[57], _091_[42], _091_[31], _091_[22], _091_[0] } = { _087_[131:123], _035_, _087_[121:0], _016_, _085_, _062_, _007_, _003_ };
  assign { _092_[34], _092_[16] } = { _068_, _028_ };
  assign { _093_[46], _093_[42], _093_[37], _093_[8] } = { _053_, _061_, _013_, _082_ };
  assign _094_[13:12] = { _046_, _026_ };
  assign { _096_[38], _096_[5:0] } = { _063_, _079_, _022_, _003_, _058_, _055_, _022_ };
  assign { _097_[46], _097_[21:0] } = { _001_, _096_[74:53] };
  assign _098_[57] = _029_;
  assign { _099_[90:27], _099_[3] } = { _095_[63:0], _059_ };
  assign _100_[128] = _057_;
  assign { _101_[168], _101_[157:0] } = { _076_, _091_[234:218], _098_[90:58], _029_, _098_[56:0], _058_, _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _079_ };
  assign _102_[32] = _021_;
  assign _104_[135:0] = { _083_, _036_, _087_[131:123], _035_, _087_[121:0], _009_, _036_ };
  assign { _105_[228:87], _105_[83], _105_[78], _105_[75:0] } = { _101_[202:169], _076_, _101_[167:158], _091_[234:204], _091_[65:58], _016_, _091_[56:43], _085_, _091_[41:32], _062_, _091_[30:23], _007_, _091_[21:1], _020_, _044_, _071_, _078_, _094_[74:14], _046_, _026_, _094_[11:0] };
  assign _106_[41] = _065_;
  assign { _107_[147:17], _107_[0] } = { _088_[131:45], _019_, _088_[43:1], _014_ };
  assign { _108_[22], _108_[19] } = { _041_, _043_ };
  assign { _109_[14], _109_[6], _109_[3:0] } = { _038_, _080_, _069_, _055_, _003_, _022_ };
  assign _110_[162] = _047_;
  assign _112_[215:0] = { _095_, _099_[26:22], _090_[174:105], _066_, _090_[103:40], _000_ };
  assign { _115_[5], _115_[1:0] } = { _031_, _069_, _011_ };
  assign { _116_[36], _116_[14] } = { _050_, _073_ };
  assign { _117_[228:25], _117_[1:0] } = { _090_[38:30], _008_, _090_[28:9], _002_, _090_[7:0], _000_, _047_, _110_[161:0], _005_, _003_, _022_ };
  assign { _119_[254], _119_[24:0] } = { _081_, _108_[23], _041_, _108_[21:20], _043_, _108_[18:0], _058_ };
  assign _120_[257:0] = { _119_[282:255], _081_, _119_[253:25] };
  assign _121_[72] = _064_;
  assign { _123_[260:224], _123_[128:126], _123_[108:16] } = { _115_[38:6], _031_, _115_[4:2], _051_, _045_, _052_, _104_[228:136] };
  assign { _124_[267:129], _124_[91:0] } = { _112_[252:216], _095_, _099_[26:4], _059_, _099_[2:0], _017_, _098_[90:58], _029_, _098_[56:0] };
  assign { _127_[219:188], _127_[156], _127_[154] } = { out_data[831:800], _060_, _067_ };
  assign _128_[202:171] = out_data[735:704];
  assign _129_[43:12] = out_data[671:640];
  assign { _130_[135:104], _130_[30] } = { out_data[639:608], _072_ };
  assign { _131_[91], _131_[81:50] } = { _077_, out_data[543:512] };
  assign { _132_[209], _132_[158:5] } = { _084_, _115_[60:6], _031_, _115_[4:2], _123_[223:129] };
  assign { _133_[124:93], _133_[58] } = { out_data[479:448], _075_ };
  assign { _134_[210:156], _134_[130:36], _134_[22], _134_[0] } = { _093_[13:10], _058_, _012_, _058_, _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], _097_[47], _001_, _097_[45:22], _096_[74:39], _063_, _096_[37:6], _010_, _012_ };
  assign { _135_[180:149], _135_[70] } = { out_data[415:384], _070_ };
  assign _136_[224:193] = out_data[383:352];
  assign _137_[38:7] = out_data[319:288];
  assign { _138_[161:58], _138_[48:0] } = { _095_[39:0], _099_[26:4], _059_, _099_[2:0], _124_[128:92], _093_[47], _053_, _093_[45:43], _061_, _093_[41:38], _013_, _093_[36:9], _082_, _093_[7:0], out_data[320] };
  assign _139_[48:17] = out_data[223:192];
  assign _140_[46:0] = { _101_[269:224], _045_ };
  assign _141_[36:5] = out_data[191:160];
  assign { _142_[278:254], _142_[246:77] } = { _087_[126:123], _035_, _087_[121:102], _107_[170:148], _088_[131:45], _019_, _088_[43:1], _107_[16:1] };
  assign _143_[162:131] = out_data[159:128];
  assign { _144_[21], _144_[19:0] } = { _040_, _109_[23:15], _038_, _109_[13:7], _080_, _109_[5:4] };
  assign _145_[249:41] = { _112_[276:216], _095_, _099_[26:4], _059_, _099_[2:0], _124_[128:92], _138_[57:49] };
  assign _146_[188:27] = { _140_[59:47], _101_[269:169], _076_, _101_[167:158], _091_[234:198] };
endmodule
